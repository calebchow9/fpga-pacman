module map_mask(
	input [8:0] x,
	input [8:0] y,
	
	output mask
);

	// ROM definition
	parameter bit [299:0] ROM [327:0]= '{
	300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000001111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
300'b 111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 };

logic [299:0] line;

assign line = ROM[y];

assign mask = line[x];

endmodule