module map_mask(
	input [9:0] x,
	input [9:0] y,
	
	output mask, 
	output [4:0] maskL, maskR, maskT, maskB
);
	logic [404:0] line;

	// maze size 405 (width) x 448 (height)
	// ROM definition
	parameter bit [404:0] bit_map [0:447]= '{
405'b 000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
405'b 000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000,
405'b 001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100,
405'b 011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111,
405'b 110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000111000000000000000000000000000000001110000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000011100000000000000000000000000000000111000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000011100000000000000000000000000000000000011100000000000000000000000000000011100000000000000000000000000000000000000000000000000011100000000000000000000000000000110000000000011000000000000000000000000000001110000000000000000000000000000000000000000000000000001110000000000000000000000000000001110000000000000000000000000000000000001110000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111100000000000000000000000000000000000011100000000000000000000000000000011100000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000001110000000000000000000000000000001110000000000000000000000000000000000001111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000111000000000000000000000000000000001110000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000011100000000000000000000000000000000111000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000011111111000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111110000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000111000000000000000000000000000000001110000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000011100000000000000000000000000000000111000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111100000000000000000000000000000000000011100000000000000000000000000000011100000001111000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000111100000001110000000000000000000000000000001110000000000000000000000000000000000001111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000011000000000000000000000000000000111000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000111000000000000000000000000000000110000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000111000000000011000000000000000000000000000000011111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111110000000000000000000000000000000110000000000111000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000111000000000011000000000000000000000000000000001111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111100000000000000000000000000000000110000000000111000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000111000000000011000000000000000000000000000000000111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111000000000000000000000000000000000110000000000111000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011110000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000011110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011,
405'b 110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000110000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011,
405'b 111100001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111000000000000111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111000000000000111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100001111,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111000000000000011111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111110000000000000111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 011100000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000111000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000111000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000001110,
405'b 001100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000111000000000000000000000000000000000000000000000000000011000000000000000000000000000000110000000000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000111000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000001100,
405'b 000111100000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000001111000,
405'b 000011111111111111111111111111111111111111111111111111111111111111111111000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000111111111111111111111111111111111111111111111111111111111111111111110000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111100001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100001111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111110001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100011111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000011000000000000000000000000000000011100000001110000000000000000000000000000000110000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000111000000000000000000000000000000001110000011100000000000000000000000000000000111000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000001111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000000001111111111111111111111111111111111111100000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000110000000000000000000000000000011000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000110000000000000000000000000000011000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000110000000000000000000000000000011000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100011111111111111111111111111111110000000000000000000000000000011111111111111111111111111111110001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000001110001110000000000000000000000000000111000000000011000000000000000000000000000001100011111111111111111111111111111110000000000000000000000000000011111111111111111111111111111110001100000000000000000000000000000110000000000111000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111100001110000000000000000000000000000111000000000011000000000000000000000000000001100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001100000000000000000000000000000110000000000111000000000000000000000000000011100001111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111000001110000000000000000000000000000111000000000011000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000110000000000111000000000000000000000000000011100000111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001111000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000111100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000001110000001100000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000001100000011100000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111100000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000001111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111111000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111111000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001110000001100000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000001100000011100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001111000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000111100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111000001110000000000000000000000000000111000000000011000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000110000000000111000000000000000000000000000011100000111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111100001110000000000000000000000000000111000000000011000000000000000000000000000001100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001100000000000000000000000000000110000000000111000000000000000000000000000011100001111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111110001110000000000000000000000000000111000000000011000000000000000000000000000001100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001100000000000000000000000000000110000000000111000000000000000000000000000011100011111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111110001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100011111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111100001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100001111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000011111111111111111111111111111111111111111111111111111111111111111111000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000111111111111111111111111111111111111111111111111111111111111111111110000,
405'b 000111110000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000011111000,
405'b 001111100000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001110000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000011100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000001111100,
405'b 011100000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001110000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000011100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000001110,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 111100001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100001111,
405'b 110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011,
405'b 110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000110000000000011000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000110000000000011000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000011000000000000000000000000000000001100000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000001100000000000000000000000000000000110000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111000000000000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000000000000000000000000000011100000000000000000000000000000110000000000011000000000000000000000000000001110000000000000000000000000000000000000000000000000001111000000000000000000000000000011110000000000000000000000000000000000000111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111100000000000000000000000000000000000001110000000000000000000000000000011100000000000000000000000000000000000000000000000000011100000000000000000000000000000111100000001111000000000000000000000000000001110000000000000000000000000000000000000000000000000001110000000000000000000000000000011100000000000000000000000000000000000001111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000001110000000000000000000000000000001100000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000001100000000000000000000000000000011100000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001111111111111111111111111000000000000001110000000000000000000000000000000111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000011100000000000000111111111111111111111111100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111100000000000001110000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000011100000000000001111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000001111111111111111111111110000000000001110000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000001111100000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000011100000000000011111111111111111111111100000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000111000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000111000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000011100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001110000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110000111000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000111000011,
405'b 110000011100000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000001110000011,
405'b 110000001111111111111111111111111000000000000000000000000000000001100000000001110000000000000000000000000000000011111111000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111110000000000000000000000000000000011100000000001100000000000000000000000000000000111111111111111111111111100000011,
405'b 110000000111111111111111111111111000000000000000000000000000000001100000000001110000000000000000000000000000000111111111000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000011100000000001100000000000000000000000000000000111111111111111111111111000000011,
405'b 110000000000000000000000000000001110000000000000000000000000000001100000000001110000000000000000000000000000001110000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000011100000000000000000000000000000011100000000001100000000000000000000000000000011100000000000000000000000000000011,
405'b 110000000000000000000000000000000111000000000000000000000000000001100000000001110000000000000000000000000000011100000001111000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000111100000001110000000000000000000000000000011100000000001100000000000000000000000000000111000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011000000000000000000000000000001110000000001110000000000000000000000000000111000000000011000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000110000000000111000000000000000000000000000011100000000011100000000000000000000000000000110000000000000000000000000000000011,
405'b 110000000000000000000000000000001110000000000000000000000000000000111000000011000000000000000000000000000000111000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000111000000000000000000000000000000110000000111000000000000000000000000000000011100000000000000000000000000000011,
405'b 110000000011111111111111111111111100000000000000000000000000000000011111111111000000000000000000000000000000111000000000011000000000000000000000000000000011111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111110000000000000000000000000000000110000000000111000000000000000000000000000000111111111110000000000000000000000000000000001111111111111111111111110000000011,
405'b 110000000111111111111111111111111000000000000000000000000000000000001111111100000000000000000000000000000000111000000000011000000000000000000000000000000001111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111100000000000000000000000000000000110000000000111000000000000000000000000000000001111111100000000000000000000000000000000000111111111111111111111111000000011,
405'b 110000011111111111111111111111110000000000000000000000000000000000000111111100000000000000000000000000000000111000000000011000000000000000000000000000000000111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111000000000000000000000000000000000110000000000111000000000000000000000000000000001111111000000000000000000000000000000000000011111111111111111111111110000011,
405'b 110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011,
405'b 110001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000110000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000011000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111000000000000000000000000000000110000000000011000000000000000000000000000000111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011,
405'b 111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,
405'b 001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100,
405'b 000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000,
405'b 000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000};

logic [9:0] offL, offR, offT, offB;
logic [404:0] lineT, lineB, lineplus, lineminus, lineminus1, lineplus1;

assign offL = x-14;
assign offR = x+14;
assign offT = y-14;
assign offB = y+14;

assign line = bit_map[y];
assign lineminus = bit_map[y-8];
assign lineminus1 = bit_map[y-12];
assign lineplus = bit_map[y+8];
assign lineplus1 = bit_map[y+12];
assign lineT = bit_map[offT];
assign lineB = bit_map[offB];

assign mask = line[x];
assign maskL = {lineminus1[offL], lineminus[offL], line[offL], lineplus[offL], lineplus1[offL]};
assign maskR = {lineminus1[offR], lineminus[offR], line[offR], lineplus[offR], lineplus1[offR]};
assign maskT = {lineT[x-11], lineT[x-8], lineT[x], lineT[x+8], lineT[x+11]};
assign maskB = {lineB[x-11], lineB[x-8], lineB[x], lineB[x+8], lineB[x+11]};

endmodule