module map_mask(
	input [9:0] x, y, rgx, rgy, ogx, ogy,
	
	output mask, 
	output [4:0] maskL, maskR, maskT, maskB, RGmaskL, RGmaskR, RGmaskT, RGmaskB, OGmaskL, OGmaskR, OGmaskT, OGmaskB
);
	logic [404:0] line;
	logic [404:0] RGline;
	logic [404:0] OGline;

	// maze size 405 (width) x 448 (height)
	// ROM definition
	parameter bit [404:0] bit_map [0:447]= '{
405'b 000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
405'b 000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000,
405'b 001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100,
405'b 011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111,
405'b 110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000111000000000000000000000000000000001110000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000011100000000000000000000000000000000111000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000011100000000000000000000000000000000000011100000000000000000000000000000011100000000000000000000000000000000000000000000000000011100000000000000000000000000000110000000000011000000000000000000000000000001110000000000000000000000000000000000000000000000000001110000000000000000000000000000001110000000000000000000000000000000000001110000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111100000000000000000000000000000000000011100000000000000000000000000000011100000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000001110000000000000000000000000000001110000000000000000000000000000000000001111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000111000000000000000000000000000000001110000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000011100000000000000000000000000000000111000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000011111111000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111110000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000111000000000000000000000000000000001110000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000011100000000000000000000000000000000111000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111100000000000000000000000000000000000011100000000000000000000000000000011100000001111000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000111100000001110000000000000000000000000000001110000000000000000000000000000000000001111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000011000000000000000000000000000000111000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000111000000000000000000000000000000110000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000111000000000011000000000000000000000000000000011111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111110000000000000000000000000000000110000000000111000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000111000000000011000000000000000000000000000000001111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111100000000000000000000000000000000110000000000111000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000111000000000011000000000000000000000000000000000111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111000000000000000000000000000000000110000000000111000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011110000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000011110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011,
405'b 110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000110000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000011000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011,
405'b 111100001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111000000000000111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111000000000000111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100001111,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111000000000000011111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111110000000000000111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 011100000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000111000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000111000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000001110,
405'b 001100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000111000000000000000000000000000000000000000000000000000011000000000000000000000000000000110000000000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000111000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000001100,
405'b 000111100000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000001111000,
405'b 000011111111111111111111111111111111111111111111111111111111111111111111000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000111111111111111111111111111111111111111111111111111111111111111111110000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111100001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100001111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111110001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100011111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000011000000000000000000000000000000011100000001110000000000000000000000000000000110000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000000000000000000000000000000000000000000111000000000000000000000000000000001110000011100000000000000000000000000000000111000000000000000000000000000000000000000000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000001111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000000001111111111111111111111111111111111111100000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000110000000000000000000000000000011000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000110000000000000000000000000000011000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000110000000000000000000000000000011000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100011111111111111111111111111111110000000000000000000000000000011111111111111111111111111111110001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000001110001110000000000000000000000000000111000000000011000000000000000000000000000001100011111111111111111111111111111110000000000000000000000000000011111111111111111111111111111110001100000000000000000000000000000110000000000111000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111100001110000000000000000000000000000111000000000011000000000000000000000000000001100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001100000000000000000000000000000110000000000111000000000000000000000000000011100001111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111000001110000000000000000000000000000111000000000011000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000110000000000111000000000000000000000000000011100000111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001111000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000111100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000001110000001100000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000001100000011100000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111100000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000001111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111111000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111111000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001110000001100000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000001100000011100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001111000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000111100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111000001110000000000000000000000000000111000000000011000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000110000000000111000000000000000000000000000011100000111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111100001110000000000000000000000000000111000000000011000000000000000000000000000001100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001100000000000000000000000000000110000000000111000000000000000000000000000011100001111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 111111111111111111111111111111111111111111111111111111111111111111111111110001110000000000000000000000000000111000000000011000000000000000000000000000001100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001100000000000000000000000000000110000000000111000000000000000000000000000011100011111111111111111111111111111111111111111111111111111111111111111111111111,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100111000000000000000000000000000000000000000000000000000000000000000000000000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111110001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100011111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111100001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100001111111111111111111111111111111111111111111111111111111111111111110000000,
405'b 000011111111111111111111111111111111111111111111111111111111111111111111000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000111111111111111111111111111111111111111111111111111111111111111111110000,
405'b 000111110000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000011111000,
405'b 001111100000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001110000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000011100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000001111100,
405'b 011100000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001110000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000011100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000001110,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 111100001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100001111,
405'b 110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011,
405'b 110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000110000000000011000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000110000000000011000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000011000000000000000000000000000000001100000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000001100000000000000000000000000000000110000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111000000000000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000000000000000000000000000011100000000000000000000000000000110000000000011000000000000000000000000000001110000000000000000000000000000000000000000000000000001111000000000000000000000000000011110000000000000000000000000000000000000111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000001110000000000000000000000000000111000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000111000000000000000000000000000011100000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111100000000000000000000000000000000000001110000000000000000000000000000011100000000000000000000000000000000000000000000000000011100000000000000000000000000000111100000001111000000000000000000000000000001110000000000000000000000000000000000000000000000000001110000000000000000000000000000011100000000000000000000000000000000000001111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000001110000000000000000000000000000001100000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000001100000000000000000000000000000011100000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001111111111111111111111111000000000000001110000000000000000000000000000000111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000011100000000000000111111111111111111111111100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111100000000000001110000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000011100000000000001111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000001111111111111111111111110000000000001110000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000001111100000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000011100000000000011111111111111111111111100000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000111000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000111000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000011100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001110000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000011100011,
405'b 110000111000000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000000111000011,
405'b 110000011100000000000000000000000000000000000000000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100000000000000000000000000000000000000000000000000000001110000011,
405'b 110000001111111111111111111111111000000000000000000000000000000001100000000001110000000000000000000000000000000011111111000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111110000000000000000000000000000000011100000000001100000000000000000000000000000000111111111111111111111111100000011,
405'b 110000000111111111111111111111111000000000000000000000000000000001100000000001110000000000000000000000000000000111111111000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000011100000000001100000000000000000000000000000000111111111111111111111111000000011,
405'b 110000000000000000000000000000001110000000000000000000000000000001100000000001110000000000000000000000000000001110000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000011100000000000000000000000000000011100000000001100000000000000000000000000000011100000000000000000000000000000011,
405'b 110000000000000000000000000000000111000000000000000000000000000001100000000001110000000000000000000000000000011100000001111000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000111100000001110000000000000000000000000000011100000000001100000000000000000000000000000111000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011100000000000000000000000000001100000000001110000000000000000000000000000111000000000011000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000110000000000111000000000000000000000000000011100000000001100000000000000000000000000001110000000000000000000000000000000011,
405'b 110000000000000000000000000000000011000000000000000000000000000001110000000001110000000000000000000000000000111000000000011000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000110000000000111000000000000000000000000000011100000000011100000000000000000000000000000110000000000000000000000000000000011,
405'b 110000000000000000000000000000001110000000000000000000000000000000111000000011000000000000000000000000000000111000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000111000000000000000000000000000000110000000111000000000000000000000000000000011100000000000000000000000000000011,
405'b 110000000011111111111111111111111100000000000000000000000000000000011111111111000000000000000000000000000000111000000000011000000000000000000000000000000011111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111110000000000000000000000000000000110000000000111000000000000000000000000000000111111111110000000000000000000000000000000001111111111111111111111110000000011,
405'b 110000000111111111111111111111111000000000000000000000000000000000001111111100000000000000000000000000000000111000000000011000000000000000000000000000000001111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111100000000000000000000000000000000110000000000111000000000000000000000000000000001111111100000000000000000000000000000000000111111111111111111111111000000011,
405'b 110000011111111111111111111111110000000000000000000000000000000000000111111100000000000000000000000000000000111000000000011000000000000000000000000000000000111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111000000000000000000000000000000000110000000000111000000000000000000000000000000001111111000000000000000000000000000000000000011111111111111111111111110000011,
405'b 110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011,
405'b 110001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000110000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000011000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111100000000000000000000000000000000110000000000011000000000000000000000000000000001111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111000000000000000000000000000000110000000000011000000000000000000000000000000111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000110000000000011000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111000000000111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000011100000001110000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000001100000001100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011,
405'b 110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011,
405'b 111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110,
405'b 011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,
405'b 001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100,
405'b 000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000,
405'b 000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
405'b 000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000};

logic [9:0] offL, offR, offT, offB;
logic [404:0] lineT, lineB, lineplus, lineminus, lineminus1, lineplus1;

assign offL = x-14;
assign offR = x+14;
assign offT = y-14;
assign offB = y+14;

assign line = bit_map[y];
assign lineminus = bit_map[y-8];
assign lineminus1 = bit_map[y-12];
assign lineplus = bit_map[y+8];
assign lineplus1 = bit_map[y+12];
assign lineT = bit_map[offT];
assign lineB = bit_map[offB];

assign mask = line[x];
assign maskL = {lineminus1[offL], lineminus[offL], line[offL], lineplus[offL], lineplus1[offL]};
assign maskR = {lineminus1[offR], lineminus[offR], line[offR], lineplus[offR], lineplus1[offR]};
assign maskT = {lineT[x-11], lineT[x-8], lineT[x], lineT[x+8], lineT[x+11]};
assign maskB = {lineB[x-11], lineB[x-8], lineB[x], lineB[x+8], lineB[x+11]};

// red ghost collisions
logic [9:0] RGoffL, RGoffR, RGoffT, RGoffB;
logic [404:0] RGlineT, RGlineB, RGlineplus, RGlineminus, RGlineminus1, RGlineplus1;

assign RGoffL = rgx-14;
assign RGoffR = rgx+14;
assign RGoffT = rgy-14;
assign RGoffB = rgy+14;

assign RGline = bit_map[rgy];
assign RGlineminus = bit_map[rgy-8];
assign RGlineminus1 = bit_map[rgy-12];
assign RGlineplus = bit_map[rgy+8];
assign RGlineplus1 = bit_map[rgy+12];
assign RGlineT = bit_map[RGoffT];
assign RGlineB = bit_map[RGoffB];

assign RGmaskL = {RGlineminus1[RGoffL], RGlineminus[RGoffL], RGline[RGoffL], RGlineplus[RGoffL], RGlineplus1[RGoffL]};
assign RGmaskR = {RGlineminus1[RGoffR], RGlineminus[RGoffR], RGline[RGoffR], RGlineplus[RGoffR], RGlineplus1[RGoffR]};
assign RGmaskT = {RGlineT[rgx-11], RGlineT[rgx-8], RGlineT[rgx], RGlineT[rgx+8], RGlineT[rgx+11]};
assign RGmaskB = {RGlineB[rgx-11], RGlineB[rgx-8], RGlineB[rgx], RGlineB[rgx+8], RGlineB[rgx+11]};

// orange ghost collisions
logic [9:0] OGoffL, OGoffR, OGoffT, OGoffB;
logic [404:0] OGlineT, OGlineB, OGlineplus, OGlineminus, OGlineminus1, OGlineplus1;

assign OGoffL = ogx-14;
assign OGoffR = ogx+14;
assign OGoffT = ogy-14;
assign OGoffB = ogy+14;

assign OGline = bit_map[ogy];
assign OGlineminus = bit_map[ogy-8];
assign OGlineminus1 = bit_map[ogy-12];
assign OGlineplus = bit_map[ogy+8];
assign OGlineplus1 = bit_map[ogy+12];
assign OGlineT = bit_map[OGoffT];
assign OGlineB = bit_map[OGoffB];

assign OGmaskL = {OGlineminus1[OGoffL], OGlineminus[OGoffL], OGline[OGoffL], OGlineplus[OGoffL], OGlineplus1[OGoffL]};
assign OGmaskR = {OGlineminus1[OGoffR], OGlineminus[OGoffR], OGline[OGoffR], OGlineplus[OGoffR], OGlineplus1[OGoffR]};
assign OGmaskT = {OGlineT[ogx-11], OGlineT[ogx-8], OGlineT[ogx], OGlineT[ogx+8], OGlineT[ogx+11]};
assign OGmaskB = {OGlineB[ogx-11], OGlineB[ogx-8], OGlineB[ogx], OGlineB[ogx+8], OGlineB[ogx+11]};

endmodule